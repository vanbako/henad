`ifndef FLAGS_VH
`define FLAGS_VH

`define FLAG_Z 0
`define FLAG_N 1
`define FLAG_C 2
`define FLAG_V 3

`endif
