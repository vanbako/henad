`include "src/sizes.vh"
`include "src/opcodes.vh"

module stg_mo(
    input wire                   iw_clk,
    input wire                   iw_rst,
    input wire  [`HBIT_ADDR:0]   iw_pc,
    output wire [`HBIT_ADDR:0]   ow_pc,
    input wire  [`HBIT_DATA:0]   iw_instr,
    output wire [`HBIT_DATA:0]   ow_instr,
    input wire  [`HBIT_OPC:0]    iw_opc,
    output wire [`HBIT_OPC:0]    ow_opc,
    input wire  [`HBIT_TGT_GP:0] iw_tgt_gp,
    input wire                   iw_tgt_gp_we,
    output wire [`HBIT_TGT_GP:0] ow_tgt_gp,
    output wire                  ow_tgt_gp_we,
    input wire  [`HBIT_TGT_SR:0] iw_tgt_sr,
    input wire                   iw_tgt_sr_we,
    output wire [`HBIT_TGT_SR:0] ow_tgt_sr,
    output wire                  ow_tgt_sr_we,
    input wire  [`HBIT_TGT_AR:0] iw_tgt_ar,
    input wire                   iw_tgt_ar_we,
    output wire [`HBIT_TGT_AR:0] ow_tgt_ar,
    output wire                  ow_tgt_ar_we,
    // iw_mem_mp selects which memory port MO uses in this cycle.
    // MA set the address on the opposite port in the previous cycle, so the
    // two ports exist to let MA and MO alternate each cycle.
    //
    // 48-bit ops do NOT use both ports simultaneously. MO still accesses a
    // single port selected by iw_mem_mp, using the full 48-bit per-port
    // buses: `ow_mem_wdata[*]` for stores and `iw_mem_rdata[*]` for loads.
    // The memory (`mem.v`) packs/unpacks adjacent 24-bit words internally
    // when `ow_mem_is48[*]` is asserted for that selected port.
    input wire                   iw_mem_mp,
    output reg                   ow_mem_we [0:1],
    output reg  [`HBIT_ADDR:0]   ow_mem_wdata [0:1],  // 48-bit write bus per port
    output reg                   ow_mem_is48 [0:1],   // per-port access width: 1=48b
    input wire  [`HBIT_ADDR:0]   iw_mem_rdata [0:1],  // 48-bit read bus per port
    input wire  [`HBIT_DATA:0]   iw_result,
    output wire [`HBIT_DATA:0]   ow_result,
    input wire  [`HBIT_ADDR:0]   iw_sr_result,
    output wire [`HBIT_ADDR:0]   ow_sr_result,
    input wire  [`HBIT_ADDR:0]   iw_ar_result,
    output wire [`HBIT_ADDR:0]   ow_ar_result
);
    reg [`HBIT_DATA:0] r_result;
    reg [`HBIT_ADDR:0] r_sr_result_next;
    reg [`HBIT_ADDR:0] r_ar_result_next;
    always @(*) begin
        ow_mem_we[0] = 1'b0;
        ow_mem_we[1] = 1'b0;
        ow_mem_wdata[0] = {`SIZE_ADDR{1'b0}};
        ow_mem_wdata[1] = {`SIZE_ADDR{1'b0}};
        ow_mem_is48[0] = 1'b0;
        ow_mem_is48[1] = 1'b0;
        r_result = iw_result;
        r_sr_result_next = iw_sr_result;
        r_ar_result_next = iw_ar_result;
        case (iw_opc)
            `OPC_SRLDso: begin
                // 48-bit little-endian load from the selected port
                // Enable 48-bit read packing on both ports to tolerate the
                // MA/MO port alternation.
                ow_mem_is48[0] = 1'b1;
                ow_mem_is48[1] = 1'b1;
                r_sr_result_next = iw_mem_rdata[iw_mem_mp];
                r_result = r_sr_result_next[23:0];
            end
            `OPC_STui, `OPC_STsi: begin
                // 24-bit store to the selected port for this cycle
                ow_mem_we[iw_mem_mp] = 1'b1;
                ow_mem_wdata[iw_mem_mp] = {24'b0, iw_result};
                ow_mem_is48[iw_mem_mp] = 1'b0;
            end
            `OPC_SRSTso: begin
                // 48-bit little-endian store on the selected port
                // Use latched SR value (from previous cycle) to align with MA
                ow_mem_we[iw_mem_mp] = 1'b1;
                ow_mem_wdata[iw_mem_mp] = r_sr_result_latch;
                ow_mem_is48[iw_mem_mp] = 1'b1;
            end
        endcase
    end
    reg [`HBIT_ADDR:0]   r_pc_latch;
    reg [`HBIT_DATA:0]   r_instr_latch;
    reg [`HBIT_OPC:0]    r_opc_latch;
    reg [`HBIT_TGT_GP:0] r_tgt_gp_latch;
    reg                  r_tgt_gp_we_latch;
    reg [`HBIT_TGT_SR:0] r_tgt_sr_latch;
    reg                  r_tgt_sr_we_latch;
    reg [`HBIT_TGT_AR:0] r_tgt_ar_latch;
    reg                  r_tgt_ar_we_latch;
    reg [`HBIT_DATA:0]   r_result_latch;
    reg [`HBIT_ADDR:0]   r_sr_result_latch;
    reg [`HBIT_ADDR:0]   r_ar_result_latch;
    always @(posedge iw_clk or posedge iw_rst) begin
        if (iw_rst) begin
            r_pc_latch        <= `SIZE_ADDR'b0;
            r_instr_latch     <= `SIZE_DATA'b0;
            r_opc_latch       <= `SIZE_OPC'b0;
            r_tgt_gp_latch    <= `SIZE_TGT_GP'b0;
            r_tgt_gp_we_latch <= 1'b0;
            r_tgt_sr_latch    <= `SIZE_TGT_SR'b0;
            r_tgt_sr_we_latch <= 1'b0;
            r_tgt_ar_latch    <= `SIZE_TGT_AR'b0;
            r_tgt_ar_we_latch <= 1'b0;
            r_result_latch    <= `SIZE_DATA'b0;
            r_sr_result_latch <= `SIZE_ADDR'b0;
            r_ar_result_latch <= `SIZE_ADDR'b0;
        end
        else begin
            r_pc_latch        <= iw_pc;
            r_instr_latch     <= iw_instr;
            r_opc_latch       <= iw_opc;
            r_tgt_gp_latch    <= iw_tgt_gp;
            r_tgt_gp_we_latch <= iw_tgt_gp_we;
            r_tgt_sr_latch    <= iw_tgt_sr;
            r_tgt_sr_we_latch <= iw_tgt_sr_we;
            r_tgt_ar_latch    <= iw_tgt_ar;
            r_tgt_ar_we_latch <= iw_tgt_ar_we;
            r_result_latch    <= r_result;
            r_sr_result_latch <= r_sr_result_next;
            r_ar_result_latch <= r_ar_result_next;
        end
    end
    assign ow_pc        = r_pc_latch;
    assign ow_instr     = r_instr_latch;
    assign ow_opc       = r_opc_latch;
    assign ow_tgt_gp    = r_tgt_gp_latch;
    assign ow_tgt_gp_we = r_tgt_gp_we_latch;
    assign ow_tgt_sr    = r_tgt_sr_latch;
    assign ow_tgt_sr_we = r_tgt_sr_we_latch;
    assign ow_tgt_ar    = r_tgt_ar_latch;
    assign ow_tgt_ar_we = r_tgt_ar_we_latch;
    assign ow_result    = r_result_latch;
    assign ow_sr_result = r_sr_result_latch;
    assign ow_ar_result = r_ar_result_latch;
endmodule
