`ifndef SR_VH
`define SR_VH

`define SR_IDX_LR  4'h0
`define SR_IDX_SSP 4'h1
`define SR_IDX_FL  4'h2
`define SR_IDX_PC  4'h3

`endif