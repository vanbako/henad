`ifndef SR_VH
`define SR_VH

`define SR_IDX_LR      2'd0
`define SR_IDX_SSP     2'd1
`define SR_IDX_PSTATE  2'd2
`define SR_IDX_FL      `SR_IDX_PSTATE
`define SR_IDX_PC      2'd3

`endif
